library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity testbench is
end testbench;

architecture tb of testbench is
	-- Here, A and B are the 16 bit input binary numbers; S is the 16 bit binary output
	-- z, 'Zero Bit', = 1 when the output S is "0000000000000000" irrespective of the carry bit
	-- c is the carry bit
	-- s0 and s1 are the Selection bits
	signal A, B, S: bit_vector(15 downto 0);
	signal z, s0, s1, c: bit;

	component ALU is
		Port(  A               : in bit_vector(15 downto 0);	-- A
				 B               : in bit_vector(15 downto 0);	-- B
				 cout            : out bit;							-- c
				 Select0, Select1: in bit; 							-- s0, s1
				 Sum             : out bit_vector(15 downto 0); -- S
				 Zero            : out bit );							-- z
	end component;

	begin 
		dut_instance: ALU
		port map(A=>A, B=>B, Sum=>S, zero => z, Select0=>s1, Select1 => s0, cout => c);

	process begin
		-- S0S1 = 00 for Addition
		-- S0S1 = 10 for Subtraction
	   -- S0S1 = 01 for NAND
	   -- S0S1 = 11 for XOR
		
		S0 <= '0';
		S1 <= '0';
		A<="0100010000011010";
		B<="0010001011111010";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="0100010000011010";
		B<="0010001011111010";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="0100010000011010";
		B<="0010001011111010";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="0100010000011010";
		B<="0010001011111010";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="0111000100000111";
		B<="0101111101011101";

		wait for 5 ns;


		S0 <= '0';
		S1 <= '1';
		A<="0111000100000111";
		B<="0101111101011101";

		wait for 5 ns;


		S0 <= '1';
		S1 <= '0';
		A<="0111000100000111";
		B<="0101111101011101";

		wait for 5 ns;


		S0 <= '1';
		S1 <= '1';
		A<="0111000100000111";
		B<="0101111101011101";

		wait for 5 ns;


		S0 <= '0';
		S1 <= '0';
		A<="0110001000001111";
		B<="1111010011111100";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="0110001000001111";
		B<="1111010011111100";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="0110001000001111";
		B<="1111010011111100";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="0110001000001111";
		B<="1111010011111100";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="0000011010010111";
		B<="1110000100101010";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="0000011010010111";
		B<="1110000100101010";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="0000011010010111";
		B<="1110000100101010";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="0000011010010111";
		B<="1110000100101010";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="1010000101111011";
		B<="0010001000110101";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="1010000101111011";
		B<="0010001000110101";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="1010000101111011";
		B<="0010001000110101";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="1010000101111011";
		B<="0010001000110101";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="1101000111111010";
		B<="0101111011101000";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="1101000111111010";
		B<="0101111011101000";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="1101000111111010";
		B<="0101111011101000";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="1101000111111010";
		B<="0101111011101000";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="1100000011100000";
		B<="1101010011111101";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="1100000011100000";
		B<="1101010011111101";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="1100000011100000";
		B<="1101010011111101";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="1100000011100000";
		B<="1101010011111101";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="1000111110010001";
		B<="1000101000100111";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="1000111110010001";
		B<="1000101000100111";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="1000111110010001";
		B<="1000101000100111";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="1000111110010001";
		B<="1000101000100111";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="0000000000000000";
		B<="0000000000000000";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="0000000000000000";
		B<="0000000000000000";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="0000000000000000";
		B<="0000000000000000";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="0000000000000000";
		B<="0000000000000000";

		wait for 5 ns;


		S0 <= '0';
		S1 <= '0';
		A<="0000000000000000";
		B<="1111111111111111";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="0000000000000000";
		B<="1111111111111111";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="0000000000000000";
		B<="1111111111111111";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="0000000000000000";
		B<="1111111111111111";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="1111111111111111";
		B<="0000000000000000";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="1111111111111111";
		B<="0000000000000000";

		wait for 5 ns;
		S0 <= '1';
		S1 <= '0';
		A<="1111111111111111";
		B<="0000000000000000";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="1111111111111111";
		B<="0000000000000000";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '0';
		A<="1111111111111111";
		B<="1111111111111111";

		wait for 5 ns;

		S0 <= '0';
		S1 <= '1';
		A<="1111111111111111";
		B<="1111111111111111";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '0';
		A<="1111111111111111";
		B<="1111111111111111";

		wait for 5 ns;

		S0 <= '1';
		S1 <= '1';
		A<="1111111111111111";
		B<="1111111111111111";

		wait for 5 ns;

	end process;
end tb;